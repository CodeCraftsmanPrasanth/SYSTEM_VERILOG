class Brand;
  local string brand;
  function new(string brand);
    this.brand=brand;
    display();
  endfunction
  local function void display();
    $display("BRAND : %0s",brand);
  endfunction
endclass

module bike;
  initial begin
    Brand b;
    b=new("HERO");
    b.display();
  end
endmodule

** Error (suppressible): (vlog-8688) design.sv(18): Illegal access to local member display.
