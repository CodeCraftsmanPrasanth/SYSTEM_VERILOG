module unpackedarray3D; 
  int  array [4][3][2]; 
  initial begin 
    foreach (array[i,k,l]) begin 
      array[i][k][l]=$random; 
    end 
    $display("array = %p",array); 
  end 
endmodule

array = '{'{'{303379748, -1064739199}, '{-2071669239, -1309649309}, '{112818957, 1189058957}}, '{'{-1295874971, -1992863214}, '{15983361, 114806029}, '{992211318, 512609597}}, '{'{1993627629, 1177417612}, '{2097015289, -482925370}, '{-487095099, -720121174}}, '{'{1924134885, -1143836041}, '{-1993157102, 1206705039}, '{2033215986, -411658546}}}
