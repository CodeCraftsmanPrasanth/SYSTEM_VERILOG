module mixedarray; 
  logic [0:1][0:3] array [5][4][3]; 
  initial begin 
    foreach (array[i,k,l,m]) begin 
      array[i][k][l][m]=$random; 
    end 
    $display("array = %p",array); 
  end 
endmodule

# array = '{'{'{'{4, 1}, '{9, 3}, '{13, 13}}, '{'{5, 2}, '{1, 13}, '{6, 13}}, '{'{13, 12}, '{9, 6}, '{5, 10}}, '{'{5, 7}, '{2, 15}, '{2, 14}}}, 
            '{'{'{8, 5}, '{12, 13}, '{13, 5}}, '{'{3, 10}, '{0, 0}, '{10, 13}}, '{'{6, 3}, '{13, 3}, '{11, 5}}, '{'{2, 14}, '{13, 15}, '{3, 10}}}, 
            '{'{'{10, 12}, '{2, 10}, '{1, 8}}, '{'{8, 9}, '{11, 6}, '{6, 14}}, '{'{12, 10}, '{11, 1}, '{5, 15}}, '{'{11, 10}, '{14, 5}, '{1, 9}}}, 
            '{'{'{2, 12}, '{15, 15}, '{8, 7}}, '{'{15, 12}, '{11, 9}, '{9, 0}}, '{'{7, 1}, '{6, 12}, '{2, 8}}, '{'{7, 13}, '{2, 14}, '{13, 9}}}, 
            '{'{'{15, 3}, '{5, 8}, '{11, 9}}, '{'{15, 10}, '{8, 6}, '{14, 12}}, '{'{10, 6}, '{3, 3}, '{15, 3}}, '{'{15, 4}, '{7, 11}, '{6, 10}}}}
