module packedarray3D;
  logic [0:4][0:3][0:2][0:3] array;
  initial begin
    foreach (array[i,k,l]) begin
      array[i][k][l]=$random;
    end
    $display("array = %p",array);
  end
endmodule

array = '{'{'{4, 1, 9}, '{3, 13, 13}, '{5, 2, 1}, '{13, 6, 13}}, '{'{13, 12, 9}, '{6, 5, 10}, '{5, 7, 2}, '{15, 2, 14}}, '{'{8, 5, 12}, '{13, 13, 5}, '{3, 10, 0}, '{0, 10, 13}}, '{'{6, 3, 13}, '{3, 11, 5}, '{2, 14, 13}, '{15, 3, 10}}, '{'{10, 12, 2}, '{10, 1, 8}, '{8, 9, 11}, '{6, 6, 14}}}
