module array2;
  int fruits [] [string];
  initial begin
    fruits = new [2];
    fruits [0] = '{ "apple" : 1, "grape" : 2 };
    fruits [1] = '{ "melon" : 3, "cherry" : 4 };
    foreach (fruits[i,fruit])  $display ("fruits[%0d][%s] = %0d", i, fruit, fruits[i][fruit]);
    $display("fruits = %p",fruits);
  end
endmodule

# fruits[0][apple] = 1
# fruits[0][grape] = 2
# fruits[1][cherry] = 4
# fruits[1][melon] = 3
# fruits = '{'{"apple":1, "grape":2 }, '{"cherry":4, "melon":3 }}
