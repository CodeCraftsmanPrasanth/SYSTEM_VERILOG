module queuearray;
  int array[$][$];
  int x[][];
  int y[0:4][0:2];
  initial begin
    array='{'{$random,$random,$random},'{$random,$random,$random},'{$random,$random,$random},'{$random,$random,$random},'{$random,$random,$random}};
    $display("array = %p",array);
    $display("array size = %0d", array.size());
    x=array;
    $display("Dynamic array = %p",x);
    y=array;
    $display("Fixed array = %p",y);
     end
endmodule

array = '{'{303379748, -1064739199, -2071669239}, '{-1309649309, 112818957, 1189058957}, '{-1295874971, -1992863214, 15983361}, '{114806029, 992211318, 512609597}, '{1993627629, 1177417612, 2097015289}}
array size = 5
Dynamic array = '{'{303379748, -1064739199, -2071669239}, '{-1309649309, 112818957, 1189058957}, '{-1295874971, -1992863214, 15983361}, '{114806029, 992211318, 512609597}, '{1993627629, 1177417612, 2097015289}}
Fixed array = '{'{303379748, -1064739199, -2071669239}, '{-1309649309, 112818957, 1189058957}, '{-1295874971, -1992863214, 15983361}, '{114806029, 992211318, 512609597}, '{1993627629, 1177417612, 2097015289}}
